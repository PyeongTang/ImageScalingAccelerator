`timescale 1ns / 1ps

module tb_top();

    reg clk, rst_n;
    reg start;
    
    wire done;
    wire run;
    wire done_led;
    wire test_us_data_valid;
    wire [23:0] test_us_data;
    wire [31:0] ram_addr;
    wire [31:0] ram_dout;
    wire ram_en;
    wire [3:0] ram_wr_en;

    top dut(
        .clk(clk),
        .rst_n(rst_n),
        .start_i(start),
        .run_o(run),
        .done_o(done),
        .done_led_o(done_led),
        .ram_addr_o(ram_addr),
        .ram_dout_o(ram_dout),
        .ram_en_o(ram_en),
        .ram_wr_en_o(ram_wr_en)
    );
    
    initial begin
        clk = 0;
        forever
            #5  clk = ~clk;
    end
    
    initial begin
        rst_n = 0;
        #300    rst_n = 1;
    end
    
    initial begin
        start = 0;
        #500    start = 1;
        #10     start = 0;
    end
   
    //-----------------------------------------------------------------------
    // I recommend you to do following things.
    // 1. Store up-sampled data into buffer.
    // 2. Generate up-sampled bmp file using buffer data.
    // 3. Load up-sampled bmp file created by reference code, 
    //    and compare it with up-sampled data generated by top module 
    //-----------------------------------------------------------------------
       
    
    //-----------------------------------------------------------------------
    // check total cycles
    //-----------------------------------------------------------------------
    reg cycle_cnt_en;
    reg cycle_cnt_done;
    reg [31:0] cycle_cnt;
    reg [31:0] cycle;
    always @ (posedge clk) begin
        if (~rst_n) begin
            cycle_cnt_en <= 0;
            cycle_cnt_done <= 0; 
        end
        else begin
            if (done) begin
                cycle_cnt_en <= 0;
                cycle_cnt_done <= 1;
            end
            else if (run) begin
                cycle_cnt_en <= 1;
            end
            else begin
                cycle_cnt_en <= 0;
                cycle_cnt_done <= 0;
            end
        end
    end
    
    always @ (posedge clk) begin
        if (~rst_n) begin
            cycle_cnt <= 0;
        end
        else begin
            if (cycle_cnt_en) begin
                cycle_cnt <= cycle_cnt + 1;
            end
            else if (cycle_cnt_done) begin
                cycle <= cycle_cnt;
                cycle_cnt <= 0;
            end
        end
    end
    
    always @(*) begin
        if (cycle_cnt_done) begin
            #20;
            $display("Total cycle: %d clock", cycle);
            $stop;
        end
    end

endmodule
